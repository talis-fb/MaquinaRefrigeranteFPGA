-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 12.1 Build 243 01/31/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Dec 09 17:43:18 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY war IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        b1 : IN STD_LOGIC := '0';
        b2 : IN STD_LOGIC := '0';
        b3 : IN STD_LOGIC := '0';
        b4 : IN STD_LOGIC := '0';
        est1 : IN STD_LOGIC := '0';
        est2 : IN STD_LOGIC := '0';
        est3 : IN STD_LOGIC := '0';
        est4 : IN STD_LOGIC := '0';
        dolar : IN STD_LOGIC := '0';
        cent : IN STD_LOGIC := '0';
        finalizado : IN STD_LOGIC := '0';
        r1 : OUT STD_LOGIC;
        r2 : OUT STD_LOGIC;
        r3 : OUT STD_LOGIC;
        r4 : OUT STD_LOGIC;
        m1 : OUT STD_LOGIC;
        m2 : OUT STD_LOGIC;
        m3 : OUT STD_LOGIC;
        m4 : OUT STD_LOGIC;
        troco : OUT STD_LOGIC;
        oo : OUT STD_LOGIC;
        oi : OUT STD_LOGIC;
        io : OUT STD_LOGIC;
        ii : OUT STD_LOGIC;
		  
		  moneySeg0 : out bit_vector(6 downto 0);
		  moneySeg1 : out bit_vector(6 downto 0);
		  
		  precoSeg0 : out bit_vector(6 downto 0);
		  precoSeg1 : out bit_vector(6 downto 0);
		  
		  sell1 : out bit_vector(6 downto 0);
		  sell2 : out bit_vector(6 downto 0);
		  sell3 : out bit_vector(6 downto 0);
		  sell4 : out bit_vector(6 downto 0)
		  	   
    );
END war;

ARCHITECTURE BEHAVIOR OF war IS
    TYPE type_fstate IS (principio,start1,start2,start3,start4,r1i05,r1EndClear,r1Troco,r2i05,r2i10,r2EndClear,r2Troco,r3i05,r3i10,r3i15,r3EndClear,r3Troco,r4i05,r4i10,r4i15,r4i20,r4EndClear,r4Troco);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 
	 signal ooS: bit;
	 signal ol: bit;
	 signal lo: bit;
	 signal ll: bit;
	 signal money: bit_vector(2 downto 0);
	 signal refrigs: bit_vector(2 downto 0);
	 
	 signal vendido: bit;
	 
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='0' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,b1,b2,b3,b4,est1,est2,est3,est4,dolar,cent,finalizado)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= principio;
            r1 <= '0';
            r2 <= '0';
            r3 <= '0';
            r4 <= '0';
            m1 <= '0';
            m2 <= '0';
            m3 <= '0';
            m4 <= '0';
            troco <= '0';
            oo <= '0';
            oi <= '0';
            io <= '0';
            ii <= '0';
        ELSE
            r1 <= '0';
            r2 <= '0';
            r3 <= '0';
            r4 <= '0';
            m1 <= '0';
            m2 <= '0';
            m3 <= '0';
            m4 <= '0';
            troco <= '0';
            oo <= '0';
            oi <= '0';
            io <= '0';
            ii <= '0';
            CASE fstate IS
                WHEN principio =>
                    IF ((((((b1 = '1') AND (b2 = '0')) AND (b3 = '0')) AND (b4 = '0')) AND (est1 = '1'))) THEN
                        reg_fstate <= start1;
                    ELSIF ((((((b1 = '0') AND (b2 = '1')) AND (b3 = '0')) AND (b4 = '0')) AND (est2 = '1'))) THEN
                        reg_fstate <= start2;
                    ELSIF ((((((b1 = '0') AND (b2 = '0')) AND (b3 = '1')) AND (b4 = '0')) AND (est3 = '1'))) THEN
                        reg_fstate <= start3;
                    ELSIF ((((((b1 = '0') AND (b2 = '0')) AND (b3 = '0')) AND (b4 = '1')) AND (est4 = '1'))) THEN
                        reg_fstate <= start4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= principio;
                    END IF;
						  
						  money<="111";
						  refrigs<="111";
						  
						  vendido<='0';
						  
						  
                WHEN start1 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r1i05;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r1EndClear;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= start1;
                    END IF;

                    r1 <= '1';
						  refrigs<="000";
						  money<="111";
						  
                WHEN start2 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r2i05;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r2i10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= start2;
                    END IF;

                    r2 <= '1';
						  refrigs<="001";
						  money<="111";
						  
                WHEN start3 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r3i05;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r3i10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= start3;
                    END IF;

                    r3 <= '1';
						  refrigs<="010";
						  money<="111";
						  
                WHEN start4 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r4i05;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r4i10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= start4;
                    END IF;

                    r4 <= '1';
						  refrigs<="011";
						  money<="111";
						  
                WHEN r1i05 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r1EndClear;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r1Troco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r1i05;
                    END IF;

                    oo <= '1';
						  ooS<= '1';
						  money<="000";
						  refrigs<="000";
						  
                WHEN r1EndClear =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r1EndClear;
                    END IF;

                    m1 <= '1';
						  money<="001";
						  refrigs<="000";
						  vendido<='1';
						  
                WHEN r1Troco =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r1Troco;
                    END IF;

                    troco <= '1';

                    m1 <= '1';
						  money<="010";
						  refrigs<="000";
						  vendido<='1';
						  
                WHEN r2i05 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r2i10;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r2EndClear;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r2i05;
                    END IF;

                    oo <= '1';
						  ooS<= '1';
						  money<="000";
						  refrigs<="001";
						  
                WHEN r2i10 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r2EndClear;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r2Troco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r2i10;
                    END IF;

                    oi <= '1';
						  ol <= '1';
						  money<="001";
						  refrigs<="001";
						  
                WHEN r2EndClear =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r2EndClear;
                    END IF;

                    m2 <= '1';
						  money<="010";
						  refrigs<="001";
						  vendido<='1';
						  
                WHEN r2Troco =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r2Troco;
                    END IF;

                    troco <= '1';

                    m2 <= '1';
						  money<="011";
						  refrigs<="001";
						  vendido<='1';
						  
                WHEN r3i05 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r3i10;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r3i15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r3i05;
                    END IF;

                    oo <= '1';
						  ooS<= '1';
						  money<="000";
						  refrigs<="010";
						  
                WHEN r3i10 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r3i15;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r3EndClear;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r3i10;
                    END IF;

                    oi <= '1';
						  ol <= '1';
						  money<="001";
						  refrigs<="010";
						  
                WHEN r3i15 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r3EndClear;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r3Troco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r3i15;
                    END IF;

                    io <= '1';
						  lo <= '1';
						  money<="010";
						  refrigs<="010";
						  
                WHEN r3EndClear =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r3EndClear;
                    END IF;

                    m3 <= '1';
						  money<="011";
						  refrigs<="010";
						  vendido<='1';
						  
                WHEN r3Troco =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r3Troco;
                    END IF;

                    troco <= '1';
						  money<="100";
						  refrigs<="010";
						  vendido<='1';

                    m3 <= '1';
                WHEN r4i05 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r4i10;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r4i15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4i05;
                    END IF;

                    oo <= '1';
						  ooS<= '1';
						  money<="000";
						  refrigs<="011";
						  
                WHEN r4i10 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r4i15;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r4i20;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4i10;
                    END IF;

                    oi <= '1';
						  ol <= '1';
						  money<="001";
						  refrigs<="011";
						  
                WHEN r4i15 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r4i20;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r4EndClear;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4i15;
                    END IF;

                    io <= '1';
						  lo <= '1';
						  money<="010";
						  refrigs<="011";
						  
                WHEN r4i20 =>
                    IF (((cent = '1') AND (dolar = '0'))) THEN
                        reg_fstate <= r4EndClear;
                    ELSIF (((cent = '0') AND (dolar = '1'))) THEN
                        reg_fstate <= r4Troco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4i20;
                    END IF;

                    ii <= '1';
						  ll <= '1';
						  money<="011";
						  refrigs<="011";
						  
                WHEN r4EndClear =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4EndClear;
                    END IF;

                    m4 <= '1';
						  money<="100";
						  refrigs<="011";
						  vendido<='1';
						  
                WHEN r4Troco =>
                    IF ((finalizado = '1')) THEN
                        reg_fstate <= principio;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= r4Troco;
                    END IF;

                    troco <= '1';
						  money<="101";
						  refrigs<="011";
						  vendido<='1';

                    m4 <= '1';
                WHEN OTHERS => 
                    r1 <= 'X';
                    r2 <= 'X';
                    r3 <= 'X';
                    r4 <= 'X';
                    m1 <= 'X';
                    m2 <= 'X';
                    m3 <= 'X';
                    m4 <= 'X';
                    troco <= 'X';
                    oo <= 'X';
                    oi <= 'X';
                    io <= 'X';
                    ii <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
	
	 
	 --money(0)<= ol or ll;
	 --money(1)<= lo or ll;
	 
	 with money select
		moneySeg0<= "1000000" when "000",
		  --gfedcba
			"1111001" when "001",
			"1111001" when "010",
			"0100100" when "011",
			"0100100" when "100",
			"0110000" when "101",
			"1000000" when "111",
			"0001001" when others;

	with money select
		moneySeg1<= "0010010" when "000",
			"1000000" when "001",
			"0010010" when "010",
			"1000000" when "011",
			"0010010" when "100",
			"1000000" when "101",
			"1000000" when "111",
			"0001001" when others;
			
--------------------------------------------------
			
	with refrigs select
		precoSeg0<= "1111001" when "000",
		  --gfedcba
			"1111001" when "001",
			"0100100" when "010",
			"0100100" when "011",
			"1000000" when "111",
			"0001001" when others;

	with refrigs select
		precoSeg1<= "1000000" when "000",
			"0010010" when "001",
			"1000000" when "010",
			"0010010" when "011",
			"1000000" when "111",
			"0001001" when others;
	 
-----------------------------------------------

	with vendido select
	sell1<=  "1111111" when '0',
				"0010010" when '1',
				"1111111" when others;

	with vendido select
	sell2<=  "1111111" when '0',
				"0000110" when '1',
				"1111111" when others;
					
	with vendido select
	sell3<=  "1111111" when '0',
				"1000111" when '1',
				"1111111" when others;

	with vendido select
	sell4<=  "1111111" when '0',
				"1000111" when '1',
				"1111111" when others;

	 
	 
END BEHAVIOR;
